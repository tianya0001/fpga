library verilog;
use verilog.vl_types.all;
entity Hell_tb is
end Hell_tb;
