library verilog;
use verilog.vl_types.all;
entity mux_3to8_tb is
end mux_3to8_tb;
