library verilog;
use verilog.vl_types.all;
entity counter_ipcore_tb is
end counter_ipcore_tb;
