library verilog;
use verilog.vl_types.all;
entity BCD_counter_top_tb is
end BCD_counter_top_tb;
