library verilog;
use verilog.vl_types.all;
entity key_tb is
end key_tb;
